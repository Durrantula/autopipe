module c432 ( clock,
	  _1, _4, _8, _11, _14, _17, _21, _24, _27, _30, _34, _37, _40, _43, _47, _50, 
	  _53, _56, _60, _63, _66, _69, _73, _76, _79, _82, _86, _89, _92, _95, _99, _102, _105, 
	  _108, _112, _115, 
	  _223, _329, _370, _421, _430, _431, _432);
	input clock; 
	input _1, _4, _8, _11, _14, _17, _21, _24, _27, _30, _34, _37, _40, _43, _47, _50, 
	_53, _56, _60, _63, _66, _69, _73, _76, _79, _82, _86, _89, _92, _95, _99, _102, _105, 
	_108, _112, _115;
	output _223, _329, _370, _421, _430, _431, _432;
	reg __c432_s__1, __c432_s__4, __c432_s__8, __c432_s__11;
	wire new_n44_, new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, 
	new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, 
	new_n58_, new_n59_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_, 
	new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, 
	new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, 
	new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, 
	new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, 
	new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, 
	new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, 
	new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, 
	new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, 
	new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, 
	new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, 
	new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, 
	new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, 
	new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, 
	new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, 
	new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, 
	new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, 
	new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, 
	new_n174_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, 
	new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, 
	new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, 
	new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, 
	new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, 
	new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, 
	new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, 
	new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, 
	new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, 
	new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, 
	new_n235_, new_n236_, new_n238_, new_n239_, new_n241_, new_n242_, 
	new_n243_, new_n244_, new_n245_, new_n246_, new_n248_, new_n249_, 
	new_n250_, new_n251_;
	wire new_w00, new_w01, new_w02, new_w03;
	assign new_n44_ = ~__c432_s__1 & __c432_s__4;
	assign new_n45_ = ~__c432_s__11 & _17;
	assign new_n46_ = ~_24 & _30;
	assign new_n47_ = ~_37 & _43;
	assign new_n48_ = ~_50 & _56;
	assign new_n49_ = ~_63 & _69;
	assign new_n50_ = ~_76 & _82;
	assign new_n51_ = ~_89 & _95;
	assign new_n52_ = ~_102 & _108;
	assign new_n53_ = ~new_n44_ & ~new_n45_;
	assign new_n54_ = ~new_n46_ & new_n53_;
	assign new_n55_ = ~new_n47_ & new_n54_;
	assign new_n56_ = ~new_n48_ & new_n55_;
	assign new_n57_ = ~new_n49_ & new_n56_;
	assign new_n58_ = ~new_n50_ & new_n57_;
	assign new_n59_ = ~new_n51_ & new_n58_;
	assign _223 = new_n52_ | ~new_n59_;
	assign new_n61_ = ~new_n44_ & ~_223;
	assign new_n62_ = new_n44_ & _223;
	assign new_n63_ = ~new_n61_ & ~new_n62_;
	assign new_n64_ = __c432_s__4 & ~__c432_s__8;
	assign new_n65_ = ~new_n63_ & new_n64_;
	assign new_n66_ = ~new_n45_ & ~_223;
	assign new_n67_ = new_n45_ & _223;
	assign new_n68_ = ~new_n66_ & ~new_n67_;
	assign new_n69_ = _17 & ~_21;
	assign new_n70_ = ~new_n68_ & new_n69_;
	assign new_n71_ = ~new_n46_ & ~_223;
	assign new_n72_ = new_n46_ & _223;
	assign new_n73_ = ~new_n71_ & ~new_n72_;
	assign new_n74_ = _30 & ~_34;
	assign new_n75_ = ~new_n73_ & new_n74_;
	assign new_n76_ = ~new_n47_ & ~_223;
	assign new_n77_ = new_n47_ & _223;
	assign new_n78_ = ~new_n76_ & ~new_n77_;
	assign new_n79_ = _43 & ~_47;
	assign new_n80_ = ~new_n78_ & new_n79_;
	assign new_n81_ = ~new_n48_ & ~_223;
	assign new_n82_ = new_n48_ & _223;
	assign new_n83_ = ~new_n81_ & ~new_n82_;
	assign new_n84_ = _56 & ~_60;
	assign new_n85_ = ~new_n83_ & new_n84_;
	assign new_n86_ = ~new_n49_ & ~_223;
	assign new_n87_ = new_n49_ & _223;
	assign new_n88_ = ~new_n86_ & ~new_n87_;
	assign new_n89_ = _69 & ~_73;
	assign new_n90_ = ~new_n88_ & new_n89_;
	assign new_n91_ = ~new_n50_ & ~_223;
	assign new_n92_ = new_n50_ & _223;
	assign new_n93_ = ~new_n91_ & ~new_n92_;
	assign new_n94_ = _82 & ~_86;
	assign new_n95_ = ~new_n93_ & new_n94_;
	assign new_n96_ = ~new_n51_ & ~_223;
	assign new_n97_ = new_n51_ & _223;
	assign new_n98_ = ~new_n96_ & ~new_n97_;
	assign new_n99_ = _95 & ~_99;
	assign new_n100_ = ~new_n98_ & new_n99_;
	assign new_n101_ = ~new_n52_ & ~_223;
	assign new_n102_ = new_n52_ & _223;
	assign new_n103_ = ~new_n101_ & ~new_n102_;
	assign new_n104_ = _108 & ~_112;
	assign new_n105_ = ~new_n103_ & new_n104_;
	assign new_n106_ = ~new_n65_ & ~new_n70_;
	assign new_n107_ = ~new_n75_ & new_n106_;
	assign new_n108_ = ~new_n80_ & new_n107_;
	assign new_n109_ = ~new_n85_ & new_n108_;
	assign new_n110_ = ~new_n90_ & new_n109_;
	assign new_n111_ = ~new_n95_ & new_n110_;
	assign new_n112_ = ~new_n100_ & new_n111_;
	assign _329 = new_n105_ | ~new_n112_;
	assign new_n114_ = ~new_n65_ & ~_329;
	assign new_n115_ = new_n65_ & _329;
	assign new_n116_ = ~new_n114_ & ~new_n115_;
	assign new_n117_ = __c432_s__4 & ~_14;
	assign new_n118_ = ~new_n63_ & new_n117_;
	assign new_n119_ = ~new_n116_ & new_n118_;
	assign new_n120_ = ~new_n70_ & ~_329;
	assign new_n121_ = new_n70_ & _329;
	assign new_n122_ = ~new_n120_ & ~new_n121_;
	assign new_n123_ = _17 & ~_27;
	assign new_n124_ = ~new_n68_ & new_n123_;
	assign new_n125_ = ~new_n122_ & new_n124_;
	assign new_n126_ = ~new_n75_ & ~_329;
	assign new_n127_ = new_n75_ & _329;
	assign new_n128_ = ~new_n126_ & ~new_n127_;
	assign new_n129_ = _30 & ~_40;
	assign new_n130_ = ~new_n73_ & new_n129_;
	assign new_n131_ = ~new_n128_ & new_n130_;
	assign new_n132_ = ~new_n80_ & ~_329;
	assign new_n133_ = new_n80_ & _329;
	assign new_n134_ = ~new_n132_ & ~new_n133_;
	assign new_n135_ = _43 & ~_53;
	assign new_n136_ = ~new_n78_ & new_n135_;
	assign new_n137_ = ~new_n134_ & new_n136_;
	assign new_n138_ = ~new_n85_ & ~_329;
	assign new_n139_ = new_n85_ & _329;
	assign new_n140_ = ~new_n138_ & ~new_n139_;
	assign new_n141_ = _56 & ~_66;
	assign new_n142_ = ~new_n83_ & new_n141_;
	assign new_n143_ = ~new_n140_ & new_n142_;
	assign new_n144_ = ~new_n90_ & ~_329;
	assign new_n145_ = new_n90_ & _329;
	assign new_n146_ = ~new_n144_ & ~new_n145_;
	assign new_n147_ = _69 & ~_79;
	assign new_n148_ = ~new_n88_ & new_n147_;
	assign new_n149_ = ~new_n146_ & new_n148_;
	assign new_n150_ = ~new_n95_ & ~_329;
	assign new_n151_ = new_n95_ & _329;
	assign new_n152_ = ~new_n150_ & ~new_n151_;
	assign new_n153_ = _82 & ~_92;
	assign new_n154_ = ~new_n93_ & new_n153_;
	assign new_n155_ = ~new_n152_ & new_n154_;
	assign new_n156_ = ~new_n100_ & ~_329;
	assign new_n157_ = new_n100_ & _329;
	assign new_n158_ = ~new_n156_ & ~new_n157_;
	assign new_n159_ = _95 & ~_105;
	assign new_n160_ = ~new_n98_ & new_n159_;
	assign new_n161_ = ~new_n158_ & new_n160_;
	assign new_n162_ = ~new_n105_ & ~_329;
	assign new_n163_ = new_n105_ & _329;
	assign new_n164_ = ~new_n162_ & ~new_n163_;
	assign new_n165_ = _108 & ~_115;
	assign new_n166_ = ~new_n103_ & new_n165_;
	assign new_n167_ = ~new_n164_ & new_n166_;
	assign new_n168_ = ~new_n119_ & ~new_n125_;
	assign new_n169_ = ~new_n131_ & new_n168_;
	assign new_n170_ = ~new_n137_ & new_n169_;
	assign new_n171_ = ~new_n143_ & new_n170_;
	assign new_n172_ = ~new_n149_ & new_n171_;
	assign new_n173_ = ~new_n155_ & new_n172_;
	assign new_n174_ = ~new_n161_ & new_n173_;
	assign _370 = new_n167_ | ~new_n174_;
	assign new_n176_ = __c432_s__1 & _223;
	assign new_n177_ = __c432_s__8 & _329;
	assign new_n178_ = _14 & _370;
	assign new_n179_ = __c432_s__4 & ~new_n176_;
	assign new_n180_ = ~new_n177_ & new_n179_;
	assign new_n181_ = ~new_n178_ & new_n180_;
	assign new_n182_ = __c432_s__11 & _223;
	assign new_n183_ = _21 & _329;
	assign new_n184_ = _27 & _370;
	assign new_n185_ = ~new_n182_ & ~new_n183_;
	assign new_n186_ = ~new_n184_ & new_n185_;
	assign new_n187_ = _17 & new_n186_;
	assign new_n188_ = _24 & _223;
	assign new_n189_ = _34 & _329;
	assign new_n190_ = _40 & _370;
	assign new_n191_ = ~new_n188_ & ~new_n189_;
	assign new_n192_ = ~new_n190_ & new_n191_;
	assign new_n193_ = _30 & new_n192_;
	assign new_n194_ = _37 & _223;
	assign new_n195_ = _47 & _329;
	assign new_n196_ = _53 & _370;
	assign new_n197_ = ~new_n194_ & ~new_n195_;
	assign new_n198_ = ~new_n196_ & new_n197_;
	assign new_n199_ = _43 & new_n198_;
	assign new_n200_ = _50 & _223;
	assign new_n201_ = _60 & _329;
	assign new_n202_ = _66 & _370;
	assign new_n203_ = ~new_n200_ & ~new_n201_;
	assign new_n204_ = ~new_n202_ & new_n203_;
	assign new_n205_ = _56 & new_n204_;
	assign new_n206_ = _63 & _223;
	assign new_n207_ = _73 & _329;
	assign new_n208_ = _79 & _370;
	assign new_n209_ = ~new_n206_ & ~new_n207_;
	assign new_n210_ = ~new_n208_ & new_n209_;
	assign new_n211_ = _69 & new_n210_;
	assign new_n212_ = _76 & _223;
	assign new_n213_ = _86 & _329;
	assign new_n214_ = _92 & _370;
	assign new_n215_ = ~new_n212_ & ~new_n213_;
	assign new_n216_ = ~new_n214_ & new_n215_;
	assign new_n217_ = _82 & new_n216_;
	assign new_n218_ = _89 & _223;
	assign new_n219_ = _99 & _329;
	assign new_n220_ = _105 & _370;
	assign new_n221_ = ~new_n218_ & ~new_n219_;
	assign new_n222_ = ~new_n220_ & new_n221_;
	assign new_n223_ = _95 & new_n222_;
	assign new_n224_ = _102 & _223;
	assign new_n225_ = _112 & _329;
	assign new_n226_ = _115 & _370;
	assign new_n227_ = ~new_n224_ & ~new_n225_;
	assign new_n228_ = ~new_n226_ & new_n227_;
	assign new_n229_ = _108 & new_n228_;
	assign new_n230_ = ~new_n187_ & ~new_n193_;
	assign new_n231_ = ~new_n199_ & new_n230_;
	assign new_n232_ = ~new_n205_ & new_n231_;
	assign new_n233_ = ~new_n211_ & new_n232_;
	assign new_n234_ = ~new_n217_ & new_n233_;
	assign new_n235_ = ~new_n223_ & new_n234_;
	assign new_n236_ = ~new_n229_ & new_n235_;
	assign _421 = ~new_n181_ & ~new_n236_;
	assign new_n238_ = ~new_n193_ & new_n199_;
	assign new_n239_ = new_n230_ & ~new_n238_;
	assign _430 = new_n205_ | ~new_n239_;
	assign new_n241_ = ~new_n193_ & ~new_n199_;
	assign new_n242_ = new_n211_ & new_n241_;
	assign new_n243_ = ~new_n205_ & new_n242_;
	assign new_n244_ = ~new_n199_ & ~new_n205_;
	assign new_n245_ = new_n217_ & new_n244_;
	assign new_n246_ = new_n230_ & ~new_n243_;
	assign _431 = new_n245_ | ~new_n246_;
	assign new_n248_ = ~new_n217_ & new_n241_;
	assign new_n249_ = new_n223_ & new_n248_;
	assign new_n250_ = ~new_n187_ & ~new_n238_;
	assign new_n251_ = ~new_n243_ & new_n250_;
	assign _432 = new_n249_ | ~new_n251_;
	assign new_w00 = _1;
	assign new_w01 = _4;
	assign new_w02 = _8;
	assign new_w03 = _11;
	always @ (posedge clock) begin
		__c432_s__1 <= new_w00;
		__c432_s__4 <= new_w01;
		__c432_s__8 <= new_w02;
		__c432_s__11 <= new_w03;
	end
endmodule
